module main
import geometry

fn main() {
	b:=geometry.Box{}
	println('Hello World! ${b.string()}')
}
