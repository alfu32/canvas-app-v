module topodb






pub const mexports=['']

